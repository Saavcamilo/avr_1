----------------------------------------------------------------------------
--
--  Test Bench for AVR
--
--  This is a test bench for the AVR entity.  The test bench
--  thoroughly tests the entity by exercising it and checking the outputs.
--  Opcode instructions are loaded through an array of std_logic_vectors,
--  and the outputs are checked similarly as well.
--
--  Revision History:
--      4/4/00   Automated/Active-VHDL    Initial revision.
--      4/4/00   Glen George              Modified to add documentation and
--                                           more extensive testing.
--     11/21/05  Glen George              Updated comments and formatting.
--      9/10/17  Camilo Saavedra          Changed some stimulus and fixed bugs
----------------------------------------------------------------------------
 

library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

library opcodes;
use opcodes.opcodes.all;


entity AVR_tb is
end AVR_tb;

architecture TB_ARCHITECTURE of AVR_tb is
    -- Component declaration of the tested unit
Component AVR is
    port(
        clk     :  in     std_logic;                        -- system clock
        RST     :  in     std_logic;                         -- Reset
		DataDB  :  inout  std_logic_vector(7 downto 0);
		ProgDB  :  in     opcode_word;
		ProgAB  :  out    std_logic_vector(15 downto 0);
		DataAB  :  out    std_logic_vector(15 downto 0);
		DataWr  :  out    std_logic;
		DataRd  :  out    std_logic
		  
    );
end Component;

    -- Stimulus signals - signals mapped to the input and inout ports of tested entity    
	 signal  clk      :  std_logic;
    -- Stimulus signals - signals mapped to the input and inout ports of tested entity    signal  Clock    :  std_logic;
    signal  Reset    :  std_logic;
    signal  DataDB   :  std_logic_vector(7 downto 0);

    -- Observed signals - signals mapped to the output ports of tested entity    signal  DataRd   :  std_logic;
    signal  DataWr   :  std_logic;
    signal  DataAB   :  std_logic_vector(15 downto 0);
    signal  ProgAB   :  std_logic_vector(15 downto 0);
    --Signal used to stop clock signal generators
    signal  END_SIM  :  BOOLEAN := FALSE;
    signal  RST      :  std_logic;
    signal  Counter  :  integer := 0;
    signal  ProgDB   :  opcode_word;
	 signal  DataRd   :  std_logic;
    -- test value types
    type  byte_array    is array (natural range <>) of std_logic_vector(7 downto 0);
    type  addr_array    is array (natural range <>) of std_logic_vector(15 downto 0);
    type  prog_array    is array (natural range <>) of std_logic_vector(15 downto 0);
-- expected data bus write signal for each instruction
signal  DataRdTestVals  :  std_logic_vector(0 to 473) :=
    "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110001100011110001100011110011110010111001111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111";

-- expected data bus read signal for each instruction
signal  DataWrTestVals  :  std_logic_vector(0 to 473) :=
    "111111111111111111111111111111111111111111111111111111111111111111111111101011011110110111110011111010111101011101011111110111101111110111010111100111001110111010101011111010111101010111101011110101111110101111010111101010101111110110111110110111110011111101101111010111101011111111111111111111111111111111111111111111111111111111111101111110010001111000100111110010001111001111100011001110000011111111111111111111111111111111111111111111111111111111111111111111111111111111";

-- supplied data bus values for each instruction (for read operations)
signal  DataDBVals      :  byte_array(0 to 327) := (
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", X"0F",      
    X"F0",      X"00",      X"05",      X"05",      X"00",      
    X"F0",      "ZZZZZZZZ", "ZZZZZZZZ", X"09",      X"00",      
    X"09",      "ZZZZZZZZ", "ZZZZZZZZ", X"09",      X"09",      
    X"09",      "ZZZZZZZZ", "ZZZZZZZZ", X"03",      X"02",      
    X"01",      "ZZZZZZZZ", "ZZZZZZZZ", X"40",      X"20",      
    X"E7",      "ZZZZZZZZ", "ZZZZZZZZ", X"26",      X"22",      
    "ZZZZZZZZ", "ZZZZZZZZ", X"16",      X"02",      "ZZZZZZZZ", 
    X"19",      X"01",      X"14",      "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", X"EE",      X"DD",      X"CC",      X"BB",      
    X"AA",      "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ", 
    "ZZZZZZZZ", "ZZZZZZZZ", "ZZZZZZZZ" );

-- expected data bus output values for each instruction (only has a value on writes)
signal  DataDBTestVals  :  byte_array(0 to 327) := (
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    X"16",      "--------", X"21",      "--------", "--------", 
    X"2D",      "--------", X"19",      "--------", "--------", 
    X"26",      "--------", X"10",      "--------",      "--------", 
    X"00",      "--------", X"02",      "--------", X"14",      
    "--------", X"08",      "--------", X"04",      "--------", 
    X"02",      "--------", "--------", "--------", "--------", 
    "--------", X"01",      "--------", "--------", X"40",      
    "--------", "--------", "--------", X"42",      "--------", 
    X"FF",      "--------", X"00",      "--------", "--------", 
    X"00",      X"01",      "--------", X"00",      X"01",      
    "--------", X"00",      "--------", "--------", X"02",      
    "--------", X"01",      "--------", X"00",      "--------", 
    X"FF",      "--------", "--------", "--------", X"FF",      
    "--------", X"00",      "--------", "--------", X"01",      
    "--------", X"02",      "--------", X"03",      "--------", 
    "--------", X"40",      "--------", X"20",      "--------", 
    "--------", X"E7",      "--------", X"19",      "--------", 
    "--------", "--------", X"FF",      "--------", X"AA",      
    "--------", "--------", X"F0",      "--------", X"FF",      
    "--------", "--------", X"87",      "--------", X"C3",      
    "--------", X"E1",      "--------", X"F0",      "--------", 
    "--------", "--------", "--------", X"09",      "--------", 
    "--------", X"09",      "--------", "--------", "--------", 
    X"09",      "--------", "--------", X"09",      "--------", 
    "--------", "--------", X"09",      X"00",      "--------", 
    "--------", "--------", "--------", X"09",      "--------", 
    "--------", X"08",      "--------", "--------", X"05",      
    "--------", X"00",      "--------", "--------", X"F0",      
    "--------", X"0F",      "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", X"AA",      "--------", "--------", "--------", 
    "--------", "--------", "--------", X"BB",      X"CC",      
    "--------", X"DD",      X"EE",      X"FF",      "--------", 
    "--------", X"AA",      X"BB",      X"CC",      "--------", 
    X"DD",      X"EE",      "--------", "--------", X"AA",      
    X"BB",      "--------", X"CC",      X"DD",      X"EE",      
    "--------", "--------", X"AA",      X"BB",      "--------", 
    "--------", X"AA",      X"BB",      X"CC",      X"AA",      
    X"BB",      X"AA",      X"BB",      X"CC",      X"DD",      
    X"EE",      "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------", "--------", "--------", 
    "--------", "--------", "--------" );

-- expected data addres bus values for each instruction
signal  DataABTestVals  :  addr_array(0 to 327) := (
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    X"0000",            "----------------", X"0001",            "----------------", "----------------", 
    X"0002",            "----------------", X"0003",            "----------------", "----------------", 
    X"0004",            "----------------", X"0005",            "----------------", "----------------", 
    X"0007",            "----------------", X"0008",            "----------------", X"0009",            
    "----------------", X"000A",            "----------------", X"000B",            "----------------", 
    X"000C",            "----------------", "----------------", "----------------", "----------------", 
    "----------------", X"000D",            "----------------", "----------------", X"000E",            
    "----------------", "----------------", "----------------", X"000F",            "----------------", 
    X"0010",            "----------------", X"0011",            "----------------", "----------------", 
    X"0012",            X"0013",            "----------------", X"0014",            X"0015",            
    "----------------", X"0016",            "----------------", "----------------", X"0017",            
    "----------------", X"0018",            "----------------", X"0019",            "----------------", 
    X"001A",            "----------------", "----------------", "----------------", X"001B",            
    "----------------", X"001C",            "----------------", "----------------", X"001D",            
    "----------------", X"001E",            "----------------", X"001F",            "----------------", 
    "----------------", X"0020",            "----------------", X"0021",            "----------------", 
    "----------------", X"0022",            "----------------", X"0023",            "----------------", 
    "----------------", "----------------", X"0024",            "----------------", X"0025",            
    "----------------", "----------------", X"0026",            "----------------", X"0027",            
    "----------------", "----------------", X"0028",            "----------------", X"0029",            
    "----------------", X"002A",            "----------------", X"002B",            "----------------", 
    "----------------", "----------------", "----------------", X"002C",            "----------------", 
    "----------------", X"002D",            "----------------", "----------------", "----------------", 
    X"002E",            "----------------", "----------------", X"002F",            "----------------", 
    "----------------", "----------------", X"0030",            X"0031",            "----------------", 
    "----------------", "----------------", "----------------", X"0032",            "----------------", 
    "----------------", X"0033",            "----------------", "----------------", X"0034",            
    "----------------", X"0035",            "----------------", "----------------", X"0036",            
    "----------------", X"0037",            "----------------", "----------------", X"0037",            
    X"0036",            X"0035",            X"0034",            X"0034",            X"0035",            
    X"0036",            "----------------", "----------------", X"0030",            X"0031",            
    X"0032",            "----------------", "----------------", X"002F",            X"002E",            
    X"002D",            "----------------", "----------------", X"001F",            X"001E",            
    X"001D",            "----------------", "----------------", X"0020",            X"0021",            
    X"0022",            "----------------", "----------------", X"0004",            X"0001",            
    "----------------", "----------------", X"0000",            X"0008",            "----------------", 
    X"0003",            X"0015",            X"0009",            "----------------", "----------------", 
    "----------------", X"0038",            "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", X"0039",            X"003A",            
    "----------------", X"003D",            X"003C",            X"003B",            "----------------", 
    "----------------", X"003E",            X"003F",            X"0040",            "----------------", 
    X"0042",            X"0041",            "----------------", "----------------", X"0043",            
    X"0044",            "----------------", X"0047",            X"0046",            X"0045",            
    "----------------", "----------------", X"0048",            X"0049",            "----------------", 
    "----------------", X"004A",            X"004B",            X"004C",            X"004D",            
    X"004E",            X"FFFF",            X"FFFE",            X"FFFD",            X"FFFC",            
    X"FFFB",            X"FFFB",            X"FFFC",            X"FFFD",            X"FFFE",            
    X"FFFF",            "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------", "----------------", "----------------", 
    "----------------", "----------------", "----------------" );

signal  ProgDBVals      :  prog_array(0 to 325) := (
"1110000000000001",
"1110000000011000",
"1110000000101001",
"1110000000111010",
"1110000001001011",
"1110000001011100",
"1110000001101101",
"1110000001111110",
"1110000010001111",
"1110000010010000",
"1110000010100000",
"1110000010110000",
"1110000011001010",
"1110000011010000",
"1110000111100100",
"1110000011110000",
"0010111000001111",
"1110000011110001",
"0010111000011111",
"1110000011110010",
"0010111000101111",
"1110000011110100",
"0010111000111111",
"1110000011111000",
"0010111001001111",
"1110000111110000",
"0010111001011111",
"1110001011110000",
"0010111001101111",
"1110010011110000",
"0010111001111111",
"1110100011110000",
"0010111010001111",
"1110101011111010",
"0010111010011111",
"1110000011111000",
"0010111010101111",
"1110100011110000",
"0010111010111111",
"1110101011111010",
"0010111011001111",
"1110111111111111",
"0010111011011111",
"1110000011111111",
"0010111011101111",
"1110111111110000",
"0010111011111111",
"1110000011110000",
"1001010000001000",
"0001111100110100",
"1001001100111101",
"0001111100110100",
"1001001100111101",
"1001010000001000",
"0001111100110100",
"1001001100111101",
"0000111101010110",
"1001001101011101",
"1001010000001000",
"0000111101010110",
"1001001101011101",
"1001011000000001",
"1001001110001101",
"1001010110100011",
"0010000000000001",
"1001001000001101",
"0010000000101110",
"1001001000101101",
"0111111111101111",
"1001001111101101",
"0111000000011000",
"1001001100011001",
"1001010001000101",
"1001001001001001",
"1001010001000101",
"1001001001001001",
"1110111100001111",
"1110000000010001",
"0000111100000001",
"1001010010001000",
"0001111100000001",
"1001001100001001",
"1111101000110011",
"1111100001110000",
"1001001001111001",
"1111101000110000",
"1001010001101000",
"1111100001110001",
"1001001001111001",
"1001010111110000",
"1001001111111001",
"1001010111110000",
"1001001111111001",
"1110000000000001",
"0001011111110000",
"1001001111111001",
"1001001100001001",
"0000011111110000",
"1001001111110001",
"1001001100000001",
"0011111111111111",
"1001001111110001",
"1110000011010011",
"1001010111011010",
"1001001111010001",
"1001010111011010",
"1001001111010001",
"1001010111011010",
"1001001111010001",
"1001010111011010",
"1001001111010001",
"1110101011011010",
"1110010111000101",
"0010011111001101",
"1001001111000001",
"0010011111001100",
"1001001111000001",
"1110000011010000",
"1001010111010011",
"1001001111010001",
"1001010111010011",
"1001001111010001",
"1001010111010011",
"1001001111010001",
"1110100011010000",
"1001010111010110",
"1001001111010001",
"1001010111010110",
"1001001111010001",
"1110000111011001",
"1001010111010001",
"1001001111010001",
"1001010111010001",
"1001001111010001",
"1110101011001010",
"1110010111010101",
"0010101111011100",
"1001001111010001",
"0010101111001100",
"1001001111000001",
"1110000011010000",
"0110111111010000",
"1001001111010001",
"0110000011011111",
"1001001111010001",
"1110000011011111",
"1001010111010111",
"1001001111010001",
"1001010111010111",
"1001001111010001",
"1001010111010111",
"1001001111010001",
"1001010111010111",
"1001001111010001",
"1110000011001010",
"1110000011010000",
"1001010000001000",
"0000101111001101",
"1001001111000001",
"1001010010001000",
"0000101111001101",
"1001001111000001",
"1110000011001010",
"1001010000001000",
"0100000011000000",
"1001001111000001",
"1001010010001000",
"0100000011000000",
"1001001111000001",
"1110000011010000",
"1110000011001010",
"1001011100100001",
"1001001111000001",
"1001001111010001",
"1110000011001010",
"1110000011010001",
"1001010000001000",
"0001101111001101",
"1001001111000001",
"1001010010001000",
"0000101111001101",
"1001001111000001",
"1110011011000100",
"0101010111001111",
"1001001111000001",
"0101000011000101",
"1001001111000001",
"1110000011001111",
"1001010111000010",
"1001001111000001",
"1001010111000010",
"1001001111000001",
"1110000010110000",
"1110001110100111",
"1001000000001100",
"1001000000001110",
"1001000000001110",
"1001000000001110",
"1001000000001101",
"1001000000001101",
"1001000000001101",
"1110000011010000",
"1110001111000000",
"1001000000011001",
"1001000000011001",
"1001000000011001",
"1110000011010000",
"1110001111000000",
"1001000000101010",
"1001000000101010",
"1001000000101010",
"1110000011110000",
"1110001011100000",
"1001000000110010",
"1001000000110010",
"1001000000110010",
"1110000011110000",
"1110001011100000",
"1001000001000001",
"1001000001000001",
"1001000001000001",
"1110000011010000",
"1110000011000000",
"1000000001011100",
"1000000001011001",
"1110000011100000",
"1110000011110000",
"1000000001100000",
"1000010001100000",
"1110000011100001",
"1000000001100010",
"1001000001110000",
"0000000000010101",
"1001000001110000",
"0000000000001001",
"1110000010110000",
"1110001110101000",
"1110101000001010",
"1001001100001100",
"1001010110100011",
"1110101100011011",
"1110110000101100",
"1110110100111101",
"1110111001001110",
"1110111101011111",
"1001001100011101",
"1001001100101101",
"1110001110101110",
"1001001100111110",
"1001001101001110",
"1001001101011110",
"1110000011010000",
"1110001111001110",
"1001001100001001",
"1001001100011001",
"1001001100101001",
"1110010011000011",
"1001001100111010",
"1001001101001010",
"1110000011110000",
"1110010011100011",
"1001001100000001",
"1001001100010001",
"1110010011101000",
"1001001100100010",
"1001001100110010",
"1001001101000010",
"1110000011010000",
"1110010011000100",
"1000001100001100",
"1000001100011101",
"1110000011110000",
"1110010011100011",
"1000001100000111",
"1000011100010000",
"1000011100100001",
"1001001100000000",
"0000000001001101",
"1001001100010000",
"0000000001001110",
"1001001100001111",
"1001001100011111",
"1001001100101111",
"1001001100111111",
"1001001101001111",
"1001000000011111",
"1001000000101111",
"1001000000111111",
"1001000001001111",
"1001000001011111",
"1100000000000001",
"0000000000000000",
"1100000000000001",
"0000000000000000",
"1001010000001000",
"1111010000001000",
"0000000000000000",
"1001010010001000",
"1111010000001000",
"0000000000000000",
"1001010010001000",
"1111000000001000",
"0000000000000000",
"1001010000001000",
"1111000000001000",
"0000000000000000",
"1110101000001010",
"1110101000011010",
"1110101100101011",
"0001001100000001",
"0000000000000000",
"0001001100000010",
"0000000000000000",
"1111110100000000",
"0000000000000000",
"1111110100000001",
"0000000000000000",
"1111111100000000",
"0000000000000000",
"1111111100000001",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000");
begin

    
    -- Unit Under Test port map
    UUT : AVR        port map  (
        clk => clk, RST => RST, DataDB => DataDB, ProgDB => ProgDB,
		ProgAB => ProgAB, DataAB => DataAB, DataWr => DataWr, DataRd => DataRd
        );
    
	 clock: process
    begin
        clk <= '1';
        wait for 5 ns; -- define a clock
        clk <= '0';
        wait for 5 ns;
    end process clock;
	 counter <= to_integer(unsigned(ProgAB));
	 main: process
	 begin
	     RST <= '0';
		  wait for 11 ns;
		  RST <= '1';
		  while counter < 325 loop
            ProgDB <= ProgDBVals(counter);
            if counter > 1 then 
            wait for 1 ns;
			assert (std_match(DataDB, DataDBTestVals(counter-1))) report "DataDB " & INTEGER'IMAGE(counter-1) & " expected " & INTEGER'IMAGE(to_integer(unsigned(DataDBTestVals(counter-1)))) & " got " & INTEGER'IMAGE(to_integer(unsigned(DataDB)));
		   assert (std_match(DataAB, DataABTestVals(counter-1))) report "DataAB " & INTEGER'IMAGE(counter-1) & " expected " & INTEGER'IMAGE(to_integer(unsigned(DataABTestVals(counter-1)))) & " got " & INTEGER'IMAGE(to_integer(unsigned(DataAB)));
            end if;
         wait until counter'event;
		   end loop;
		    ProgDB <= "0000000000000000";
          wait for 10000 ns;
    end process;
end architecture;